// MOTE: This file was generated with the command:
// icepll -m -i 12 -o 30

/**
 * PLL configuration
 *
 * This Verilog module was generated automatically
 * using the icepll tool from the IceStorm project.
 * Use at your own risk.
 *
 * Given input frequency:        12.000 MHz
 * Requested output frequency:   30.000 MHz
 * Achieved output frequency:    30.000 MHz
 */

module pll (
    input  clock_in,
    output clock_out,
    output locked
);

  SB_PLL40_CORE #(
      .FEEDBACK_PATH("SIMPLE"),
      .DIVR(4'b0000),  // DIVR =  0
      .DIVF(7'b1001111),  // DIVF = 79
      .DIVQ(3'b101),  // DIVQ =  5
      .FILTER_RANGE(3'b001)  // FILTER_RANGE = 1
  ) pll_core (
      .LOCK(locked),
      .RESETB(1'b1),
      .BYPASS(1'b0),
      .REFERENCECLK(clock_in),
      .PLLOUTCORE(clock_out),

      // Unused
      .PLLOUTGLOBAL(),
      .EXTFEEDBACK(),
      .LATCHINPUTVALUE(),
      .SDO(),
      .SDI(),
      .SCLK(),
      .DYNAMICDELAY()

  );

endmodule

