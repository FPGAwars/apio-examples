module and_gate (
    input  logic a,
    input  logic b,
    output logic s
);

  assign s = a & b;

endmodule
