//--------------------------------------
//-- Turning on the LED
//--------------------------------------

module top(
    output led,   //-- LEDs
);

  // Turn on the led
  // (output the bit 1 to the led)
  assign led = 1'b1;

endmodule

