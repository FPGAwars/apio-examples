//--------------------------------------
//-- Turning on the LED
//--------------------------------------

module top(
    output led,   //-- LEDs
);

  // Turn on the led
  // (output the bit 0 to the led)
  assign led = 1'b0;

endmodule

