//------------------------------------------------------------------
//-- Verilog template
//-- Top entity
//-- Board: icezum
//------------------------------------------------------------------
`default_nettype none

//-- Template for the top entity
module top (
    output wire LED0
);

  //-- Turn on the LED0 on the icezum
  assign LED0 = 1'b1;

endmodule
