//------------------------------------------------------------------
//-- Hello world example for the EDU-CIAA-FPGA
//-- Turn on the green LED
//------------------------------------------------------------------
module leds(output wire LEDG);
 
  assign LEDG = 1'b1;
  
endmodule

