//------------------------------------------------------------------
//-- Blinking LED
//------------------------------------------------------------------

module Test (
    input  CLK,  // 25MHz clock
    output led   // LED to blink
);

  reg [23:0] counter = 0;

  always @(posedge CLK) counter <= counter + 1;

  assign led = counter[23];

endmodule
